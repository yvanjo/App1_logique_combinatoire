----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05/12/2021 12:36:34 AM
-- Design Name: 
-- Module Name: decodeur3_8_adder - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity decodeur3_8_adder is
  Port ( A : in std_logic_vector (2 downto 0);
   B : out std_logic_vector (7 downto 0));
end decodeur3_8_adder;

architecture Behavioral of decodeur3_8_adder is

begin
--process (A)
    --begin 
        --case A is
        with A select B <=
        "00000001" when "000",
        "00000010" when "001",
        "00000100"  when "010",
       "00001000" when "011" ,
        "00010000" when "100" ,
        "00100000" when "101",
        "01000000" when "110",
        "10000000"  when "111",
        "00000000" when others;

end Behavioral;
